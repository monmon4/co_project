
module SIGN_EXT (Out,In);

   input wire [15:0] In;
   output  [31:0] Out;
   
   assign Out = In;  

   
endmodule
